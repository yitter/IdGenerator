module contract

pub interface IIdGenerator {
	new_long() u64
}
