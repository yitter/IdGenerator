module contract

pub interface ISnowWorker {
	next_id() u64
}
